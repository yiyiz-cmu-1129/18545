module video_ram(
	input logic [15:0] MA;
	input logic VRAM_4HDL;
);

endmodule
