module video_ram(

);

endmodule
